always@(*) begin
    state_nxt = state;

    case(state)
    

    default: begin

    end
    endcase
end
