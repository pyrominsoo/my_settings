always@(posedge clk or negedge rstn) begin
    if (~rstn) begin

    end
    else begin

    end
end
