always@(*) begin

end
