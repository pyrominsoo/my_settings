module modulename
#(
    parameter
)
(
    input clk,
    input rstn,

);
// Registers


// Wires


endmodule
